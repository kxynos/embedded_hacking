// FPGA
// Coded by Konstantinos Xynos (2020)
// MIT License 
// Based on the blink led demo provided with Tinyfpga 
//
// look in pins.pcf for all the pin names on the TinyFPGA BX board
module out_pin (
    input CLK,    // 16MHz clock
    output PIN_1,
    output LED,   // User/boot LED next to power LED
    output USBPU  // USB pull-up resistor

);
    // drive USB pull-up resistor to '0' to disable USB
    assign USBPU = 0;

    ////////
    // make a simple blink circuit
    ////////

    // keep track of time and location in blink_pattern
    reg [25:0] blink_counter;

    // pattern that will be flashed over the LED over time
    wire [31:0] blink_pattern = 32'b101010001110111011100010101;

    // increment the blink_counter every clock
    always @(posedge CLK) begin
        blink_counter <= blink_counter + 1;
    end

    // light up the LED according to the pattern
    assign LED = blink_pattern[blink_counter[25:21]];

    // send the blink_pattern to PIN_1
    assign PIN_1 = blink_pattern[blink_counter[25:21]];
endmodule
